��     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.4.1.post1�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK
��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K
�
_n_samples�K��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�K��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��h3�f8�����R�(KhPNNNJ����J����K t�b�C              �?�t�bhTh'�scalar���hOC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���K
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hK�
node_count�K!�nodes�h)h,K ��h.��R�(KK!��h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h�h3�i8�����R�(KhPNNNJ����J����K t�bK ��h�h�K��h�h�K��h�haK��h�haK ��h�h�K(��h�haK0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@                	             �?z�):���?^            �b@                                   �?>A�F<�?/             S@                                  d@:ɨ��?            �@@                               ����?���N8�?             5@                                  �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     &@        	       
                   �i@      �?             (@        ������������������������       �                     �?                                   �D@"pc�
�?             &@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  �p@�ʈD��?            �E@                                 `c@(;L]n�?             >@       ������������������������       �                     =@        ������������������������       �                     �?                                  (q@�θ�?             *@        ������������������������       �                     @        ������������������������       �                     $@                                  �o@�����?/            �R@       ������������������������       �                      H@                                  0p@R�}e�.�?             :@        ������������������������       �                     @                                  �c@�㙢�c�?             7@        ������������������������       �                     &@                                   �?�q�q�?             (@        ������������������������       �                      @                                    d@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �t�b�values�h)h,K ��h.��R�(KK!KK��ha�B  H�z�G�?q=
ףp�?Cy�5��?������?e�M6�d�?N6�d�M�?�a�a�?��y��y�?�������?�������?              �?      �?                      �?      �?      �?              �?/�袋.�?F]t�E�?      �?      �?              �?      �?              �?        �}A_з?A_���?�?�������?              �?      �?        �؉�؉�?ى�؉��?      �?                      �?�Ϻ���?v�)�Y7�?      �?        'vb'vb�?�;�;�?              �?�7��Mo�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK!hyh)h,K ��h.��R�(KK!��h��B@                	             �?�bˢ�?d            �b@                                   �?������?2            �R@                                   n@R�}e�.�?             :@                                   �?���Q��?
             $@                                 �g@      �?              @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                     @        	       
                    �?�q�q�?             @        ������������������������       �                     �?                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                ����?      �?
             0@                                  �?      �?              @       ������������������������       �                     @                                  �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   @M@@��8��?             H@       ������������������������       �                     A@                                  `b@@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?                                   �c@�"w����?2             S@                                  @O@P�Lt�<�?             C@       ������������������������       �                    �A@                                  �t@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     C@        �t�bh�h)h,K ��h.��R�(KK!KK��ha�B  ��N��?��b�/��?к����?��g�`��?�;�;�?'vb'vb�?333333�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?      �?      �?      �?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?�$I�$I�?n۶m۶�?              �?      �?        Cy�5��?(�����?���k(�?(�����?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK1hyh)h,K ��h.��R�(KK1��h��B@                             �?�O�y���?b            �b@                      	             �?      �?             D@               
                   �j@�eP*L��?             &@                     	             �?r�q��?             @        ������������������������       �                     �?                                   a@z�G�z�?             @        ������������������������       �                      @               	                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  @e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     =@                                pff�?��̀�R�?F            �[@                      	             �?J��D��?              K@                                   _@�8��8��?             (@        ������������������������       �                     @                                  �n@؇���X�?             @                                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �J@؇���X�?             E@       ������������������������       �                     9@                                  0e@ҳ�wY;�?	             1@       ������������������������       �                     $@                                   �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?               (                    @K@�>4և��?&             L@                #                    �?�ՙ/�?             5@        !       "                   �^@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        $       %                    @I@؇���X�?             ,@       ������������������������       �                     "@        &       '                    �I@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        )       *                 ����? >�֕�?            �A@       ������������������������       �                     0@        +       ,                    a@�KM�]�?
             3@        ������������������������       �                     (@        -       0                    @N@����X�?             @        .       /                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK1KK��ha�B  ~��K~�?�6�i�?      �?      �?t�E]t�?]t�E�?�������?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?              �?        X���oX�?T�<%�S�?�^B{	��?_B{	�%�?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?        �$I�$I�?۶m۶m�?              �?      �?        �m۶m��?�$I�$I�?�a�a�?�<��<��?۶m۶m�?�$I�$I�?              �?      �?        �$I�$I�?۶m۶m�?              �?�������?333333�?      �?                      �?�A�A�?��+��+�?              �?(�����?�k(���?              �?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK-hyh)h,K ��h.��R�(KK-��h��B@                             �?� �	��?`            �b@                     	             �?�ĚpF�?9            @U@                                   \@�>4և��?             <@        ������������������������       �                     &@                                   `@�t����?             1@        ������������������������       �                      @                                ����?z�G�z�?	             .@                                  �y@      �?              @       	       
                    b@���Q��?             @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?x�}b~|�?)            �L@                                   a@      �?             @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                   �O@`'�J�?%            �I@       ������������������������       �        #             H@                                   c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               ,                    @��ɉ�?'            @P@              !                 ����?      �?&             P@                                   @J@�eP*L��?             &@        ������������������������       �                     @                       	             �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        "       )                    �?�&=�w��?!            �J@       #       $                   �p@@�E�x�?            �H@       ������������������������       �                     A@        %       &                   @a@��S�ۿ?	             .@       ������������������������       �                     "@        '       (                   �q@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        *       +                   �h@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK-KK��ha�B�  )\���(�?�Q����?uuuuuu�?�?�m۶m��?�$I�$I�?              �?�������?�������?      �?        �������?�������?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�YLg1�?Lg1��t�?      �?      �?      �?      �?      �?                      �?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�����?�����?      �?      �?t�E]t�?]t�E�?              �?۶m۶m�?�$I�$I�?              �?      �?        �x+�R�?tHM0���?9/���?և���X�?              �?�?�������?              �?UUUUUU�?�������?      �?                      �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hK
hxK-hyh)h,K ��h.��R�(KK-��h��B@                	             �?�EH,���?_            �b@                                   �R@h�˹�?+             S@                                   C@�����?*            �R@        ������������������������       �                     �?                                  �c@�F��O�?)            @R@                                 �k@�i�y�?#            �O@        ������������������������       �                     9@                                   �?�}�+r��?             C@        	                            O@����X�?             @       
                           �J@r�q��?             @                                 �_@�q�q�?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ?@                                  `d@���Q��?             $@                                   �?      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               ,                    @��(�2Y�?4            �R@              #                    �?���Hx�?3             R@                                   �n@����X�?
             ,@        ������������������������       �                     @        !       "                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        $       %                    @M@�8���?)             M@       ������������������������       �        #            �H@        &       '                   Pc@�q�q�?             "@        ������������������������       �                     @        (       +                   �q@      �?             @       )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK-KK��ha�B�  �_,�Œ�?7�i�6�?�5��P�?^Cy�5�?v�)�Y7�?�Ϻ���?      �?        �P�B�
�?�իW�^�?AA�?�������?              �?(�����?�5��P�?�$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?      �?                      �?�������?333333�?      �?      �?      �?      �?              �?      �?              �?        UUUUUU�?�������?              �?      �?              �?        �����?*�Y7�"�?9��8���?9��8��?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?j��FX�?a���{�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxKhyh)h,K ��h.��R�(KK��h��B�                	             �?�bˢ�?^            �b@                                  �c@�ӭ�a��?*             R@                                  �?P���Q�?#             N@       ������������������������       �                    �I@                                   �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @                                   �?�q�q�?             (@       	                          pe@���Q��?             $@        
                          �^@�q�q�?             @        ������������������������       �                      @                      	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                   �?$�q-�?4            �S@                                833@�����?             3@                                 `c@     ��?
             0@                                  �H@@4և���?             ,@                                  �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        )            �M@        �t�bh�h)h,K ��h.��R�(KKKK��ha�B�  ��N��?��b�/��?�8��8��?�q�q�?�������?ffffff�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?        �؉�؉�?;�;��?Q^Cy��?^Cy�5�?      �?      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK%hyh)h,K ��h.��R�(KK%��h��B@	                             �?�X�Ĳ��?_            �b@                                  �?�������?<            �V@                                  �_@*;L]n�?             >@        ������������������������       �                     $@                      	             �?��Q��?             4@                                  `@�<ݚ�?             "@        ������������������������       �                     �?                                    G@      �?              @        	       
                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@                                   �M@��S�ۿ?*             N@                                  �J@�O4R���?$            �J@       ������������������������       �                    �D@                                   g@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?                                   �?և���X�?             @        ������������������������       �                     @                                  �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                ����?r�q��?#             N@                                   @K@�<ݚ�?             "@        ������������������������       �                     �?                                  p@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                    c@�IєX�?            �I@       ������������������������       �                    �E@        !       $                    @      �?              @       "       #                    d@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK%KK��ha�BP  �@�t��?K~��K�?�������?�������?�������?""""""�?              �?�������?ffffff�?�q�q�?9��8���?      �?              �?      �?      �?      �?              �?      �?                      �?      �?        �������?�?:�&oe�?�x+�R�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?UUUUUU�?�������?9��8���?�q�q�?              �?      �?      �?              �?      �?        �?�?              �?      �?      �?333333�?�������?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK'hyh)h,K ��h.��R�(KK'��h��B�	                 	             �?�EH,���?e            �b@              	                    �?r�q��?7             U@                                   �?j���� �?	             1@                                  �g@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        
                           �?pH����?.            �P@                                  Pa@�d�����?             3@                                 �`@�q�q�?             .@                                   O@����X�?             ,@                                 �\@"pc�
�?             &@                                  �r@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   @M@ �q�q�?             H@       ������������������������       �                     ?@                      	             �?�t����?
             1@        ������������������������       �                     @                                  �n@z�G�z�?             $@       ������������������������       �                     @                                  �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        !       "                    �L@�C��2(�?.            �P@       ������������������������       �        $            �I@        #       &                    �M@���Q��?
             .@        $       %                   hu@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK'KK��ha�Bp  �_,�Œ�?7�i�6�?UUUUUU�?�������?ZZZZZZ�?�������?۶m۶m�?�$I�$I�?              �?      �?        �������?�������?              �?      �?        z�rv��?�1���?y�5���?Cy�5��?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?UUUUUU�?�������?              �?�?<<<<<<�?              �?�������?�������?              �?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?        333333�?�������?�$I�$I�?۶m۶m�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK1hyh)h,K ��h.��R�(KK1��h��B@                             �?��S���?[            �b@                                 t@�I� �?8             W@              
       	             �?���� �?3            �T@                                   �?�����H�?             2@        ������������������������       �                     @               	                   �e@"pc�
�?             &@                                  @O@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?                                pff�?     ��?'             P@                                 �f@@3����?"             K@       ������������������������       �        !            �J@        ������������������������       �                     �?                                   �?      �?             $@        ������������������������       �                     @                                ����?r�q��?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  @_@z�G�z�?             $@                                  ({@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     @               0                   �u@\-��p�?#             M@              )                 033�?���5��?"            �L@               "                    k@�θ�?             :@                !                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        #       (                    c@�KM�]�?             3@       $       %                    �M@�X�<ݺ?
             2@       ������������������������       �                     .@        &       '                    �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        *       +                   �p@�g�y��?             ?@       ������������������������       �                     9@        ,       -                 ����?r�q��?             @        ������������������������       �                     @        .       /                   s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK1KK��ha�B  �������?�?Y�B���?Nozӛ��?jW�v%j�?,Q��+�?�q�q�?�q�q�?              �?F]t�E�?/�袋.�?�������?�������?              �?      �?              �?              �?      �?���Kh�?h/�����?      �?                      �?      �?      �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?                      �?      �?      �?      �?                      �?�{a���?a����?��Gp�?�}��?�؉�؉�?ى�؉��?�$I�$I�?۶m۶m�?      �?                      �?(�����?�k(���?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �B!��?��{���?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK)hyh)h,K ��h.��R�(KK)��h��B@
                	             �?�bˢ�?`            �b@               	                    �?>A�F<�?0             S@                                  �m@���|���?             &@                                 �g@      �?              @                                  �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        
                          �\@ ����?)            @P@                                  �e@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @                                   �?�NW���?#            �J@                                  ``@     ��?             0@       ������������������������       �                     &@                                  �`@���Q��?             @        ������������������������       �                      @                                @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   c@�?�|�?            �B@       ������������������������       �                     A@                                  Pc@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?,N�_� �?0            �R@        ������������������������       �                     ;@               $                    �?�*/�8V�?            �G@                                  ``@�	j*D�?             *@        ������������������������       �                     @                #                 833@      �?              @       !       "                   `e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        %       &                     M@г�wY;�?             A@       ������������������������       �                     ?@        '       (                   0`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK)KK��ha�B�  ��N��?��b�/��?Cy�5��?������?]t�E]�?F]t�E�?      �?      �?      �?      �?      �?                      �?      �?                      �?�����?�ȍ�ȍ�?      �?      �?              �?      �?        �x+�R�?萚`���?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?к����?*�Y7�"�?              �?UUUUUU�?UUUUUU�?      �?                      �?h�`�|��?���L�?      �?        r1����?m�w6�;�?vb'vb'�?;�;��?      �?              �?      �?�������?�������?      �?                      �?              �?�?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxKhyh)h,K ��h.��R�(KK��h��B@                          `ff�?v�(��O�?]            �b@                                   Q@l{��b��?3            �S@                     	             �? ��Ou��?2            �S@                                  `m@���Q��?             $@                                 �g@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        	       
                   �r@ ��ʻ��?+             Q@       ������������������������       �        #             L@                                   �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?                                   �?O�o9%�?*            �Q@       ������������������������       �                    �I@                                pff�?��Q��?             4@                     	             �?؇���X�?             ,@                                  �c@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKKK��ha�B�  Y�%�X�?O贁N�?${�ґ�?�&��jq�?.��-���?�i�i�?333333�?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��RO�o�?�D+l$�?              �?�������?ffffff�?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?              �?      �?              �?        UUUUUU�?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK!hyh)h,K ��h.��R�(KK!��h��B@                             �?�X�Ĳ��?]            �b@                               pff�?�՘���?<            �W@              
                    �?PN��T'�?4            @T@                                  �_@p�ݯ��?             3@        ������������������������       �                     @               	                   �_@؇���X�?
             ,@                                  `c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@                                   �?6uH���?'             O@                                   `@      �?             @        ������������������������       �                      @                                   d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �c@XB���?$             M@       ������������������������       �        !             I@                                   �?      �?              @       ������������������������       �                     @        ������������������������       �                      @                                   �K@����X�?             ,@                      	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                    @lGts��?!            �K@                     	             �?�NW���?             �J@       ������������������������       �                     G@                                   @I@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK!KK��ha�B  �@�t��?K~��K�?n�S���?Fڱa��?&���^B�?h/�����?^Cy�5�?Cy�5��?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        k���Zk�?��RJ)��?      �?      �?              �?      �?      �?      �?                      �?GX�i���?�{a���?      �?              �?      �?      �?                      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?�־a�?�<%�S��?�x+�R�?萚`���?              �?�$I�$I�?۶m۶m�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hK
hxK=hyh)h,K ��h.��R�(KK=��h��B@                             @K@      �?d            �b@                                 Pm@=&C��?9            �T@              
                 433�?��<b���?             G@              	       	             �?�FVQ&�?            �@@                                  0e@      �?             @        ������������������������       �                     �?                                  pe@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@                                   �?�n_Y�K�?
             *@       ������������������������       �                     @                                033�?r�q��?             @                                   �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?��+��?            �B@                                  �?      �?             8@        ������������������������       �                      @                      	             �?"pc�
�?             6@                                  �e@      �?              @                                 ``@z�G�z�?             @        ������������������������       �                      @                                  �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �        	             *@               <                   (u@�%o��?+            �P@               3                 `ff�?     ��?)             P@        !       2                   �d@���>4��?             <@       "       1                    @8�A�0��?             6@       #       ,       	             �?�\��N��?             3@        $       +                    �?���!pc�?             &@       %       &                 ����?���Q��?             @        ������������������������       �                     �?        '       *                     O@      �?             @       (       )                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        -       .                   �`@      �?              @        ������������������������       �                     @        /       0                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        4       5                    �?�8��8��?             B@       ������������������������       �                     >@        6       7                    �O@      �?             @        ������������������������       �                      @        8       9                    �Q@      �?             @        ������������������������       �                      @        :       ;                 033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK=KK��ha�B�        �?      �?�%���?�����\�?��,d!�?��Moz��?>����?|���?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ى�؉��?;�;��?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?        *�Y7�"�?�S�n�?      �?      �?              �?/�袋.�?F]t�E�?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?\�՘H�?���[��?      �?      �?I�$I�$�?n۶m۶�?/�袋.�?颋.���?�5��P�?y�5���?t�E]t�?F]t�E�?333333�?�������?              �?      �?      �?      �?      �?              �?      �?              �?                      �?      �?      �?      �?        333333�?�������?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK/hyh)h,K ��h.��R�(KK/��h��B�                	             �?�bˢ�?a            �b@                                  �c@l{��b��?0            �S@              
                    c@��?^�k�?(            �Q@                                  �?     ��?$             P@       ������������������������       �                     H@               	                    �?      �?
             0@                                ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@                      	             �?r�q��?             @        ������������������������       �                     @                                  �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   @N@X�<ݚ�?             "@                                 �`@�q�q�?             @                                  �\@�q�q�?             @        ������������������������       �                     �?                                  �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               .                   �g@D��\��?1            �Q@              %                    �?ДX��?0             Q@               "                    �L@�t����?             1@                                  �?8�Z$���?
             *@       ������������������������       �                     "@                                  �l@      �?             @        ������������������������       �                     �?                !                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #       $                   �`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        &       -                    @`'�J�?$            �I@       '       (                    d@p���?#             I@       ������������������������       �                     A@        )       ,                   Pd@      �?             0@        *       +                     L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK/KK��ha�B�  ��b�/��?��N��?�&��jq�?${�ґ�?�A�A�?_�_��?      �?     ��?              �?      �?      �?      �?      �?      �?                      �?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?�o�z2~�?�@�6�?�������?ZZZZZZ�?�������?�������?;�;��?;�;��?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �������?�?\���(\�?{�G�z�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK+hyh)h,K ��h.��R�(KK+��h��B�
         "                 033�?Fx$(�?_            �b@                     	             �?��<b���?G            �\@               
                    �?��
P��?            �A@                               ����?���|���?             6@                                   F@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @               	                   �b@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?                                  �c@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @                                   �L@p=
ףp�?4             T@                                  �?0�z��?�?)             O@       ������������������������       �        $            �K@                                  ``@؇���X�?             @                               @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  �i@�q�q�?             2@        ������������������������       �                      @                                   �?      �?
             0@        ������������������������       �                     @               !                   �b@���Q��?             $@                                  �?�q�q�?             "@                                @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        #       &                    �?�#-���?            �A@        $       %                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        '       (                   `b@XB���?             =@       ������������������������       �                     ;@        )       *                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK+KK��ha�B�  ףp=
��?R���Q�?��,d!�?��Moz��?_�_��?PuPu�?]t�E]�?F]t�E�?333333�?ffffff�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?ى�؉��?              �?      �?        333333�?ffffff�?|���{�?�B!��?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        333333�?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?                      �?              �?_�_�?�A�A�?UUUUUU�?UUUUUU�?      �?                      �?�{a���?GX�i���?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK;hyh)h,K ��h.��R�(KK;��h��B�         *                    �?X���[�?_            �b@                                  �?�3Ea�$�?>             W@                                ����?h+�v:�?             A@                                 �|@      �?             <@                     	             �?�<ݚ�?             ;@                                   �?�n_Y�K�?             *@        ������������������������       �                     @               	                    �?z�G�z�?             $@        ������������������������       �                     �?        
                           �M@�����H�?             "@       ������������������������       �                     @                                  �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �d@@4և���?             ,@       ������������������������       �        
             *@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               '                   �g@��ϭ�*�?'             M@              &                 ���@@4և���?%             L@              #                    @�1�`jg�?$            �K@                                  �? ��WV�?!             J@        ������������������������       �                     =@                                  @a@���}<S�?             7@       ������������������������       �        
             0@               "                 ����?����X�?             @              !                   d@���Q��?             @                     	             �?�q�q�?             @        ������������������������       �                     �?                                   `a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        $       %                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        (       )                   pn@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        +       :                   �c@8^s]e�?!             M@       ,       9                    @Jm_!'1�?            �H@       -       2                    @M@�C��2(�?             F@       .       1                 ����?�g�y��?             ?@        /       0                    �I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     <@        3       6                    �M@�θ�?             *@        4       5                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       8                   �s@ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KK;KK��ha�B�  ��:m��?�X�%��?����7��?��,d!�?�������?xxxxxx�?      �?      �?9��8���?�q�q�?;�;��?ى�؉��?              �?�������?�������?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        n۶m۶�?�$I�$I�?      �?                      �?              �?              �?����=�?|a���?n۶m۶�?�$I�$I�?A��)A�?�־a�?O��N���?;�;��?      �?        ӛ���7�?d!Y�B�?      �?        �m۶m��?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?	�=����?|a���?������?����X�?F]t�E�?]t�E�?�B!��?��{���?UUUUUU�?UUUUUU�?              �?      �?                      �?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK-hyh)h,K ��h.��R�(KK-��h��B@                             �?      �?e            �b@                                 �Z@�d�����??            �W@                                   g@      �?              @                                  �W@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                      	             �?V�a�� �?:            �U@        	                          pe@8�A�0��?             6@       
                          �g@�����?             3@        ������������������������       �                     @                                  Po@և���X�?	             ,@                                 0e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �\@      �?              @        ������������������������       �                     @                                  �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   f@$�q-�?,            @P@                                  �L@���N8�?+            �O@       ������������������������       �        $            �I@                                   �?      �?             (@        ������������������������       �                      @                                   �P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               *                   �u@�C��2(�?&            �K@               '       	             �?`2U0*��?$             I@       !       "                    @M@@��8��?"             H@       ������������������������       �                     :@        #       $                   b@���7�?             6@       ������������������������       �                     4@        %       &                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        +       ,       	             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK-KK��ha�B�        �?      �?Cy�5��?y�5���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?��{a�?a���{�?/�袋.�?颋.���?^Cy�5�?Q^Cy��?              �?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?      �?              �?      �?      �?      �?                      �?      �?        �؉�؉�?;�;��?��y��y�?�a�a�?      �?              �?      �?      �?              �?      �?              �?      �?                      �?F]t�E�?]t�E�?{�G�z�?���Q��?UUUUUU�?UUUUUU�?              �?F]t�E�?�.�袋�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?        333333�?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK3hyh)h,K ��h.��R�(KK3��h��B�                	             �?*!�,��?Y            �b@                                   �B@�A+K&:�?,             S@                                  �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?z��R[�?*            �Q@                                  c@X�;�^o�?             �K@                                  �?`Ql�R�?            �G@        	                           �?z�G�z�?             @       
                          �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     E@                                `ff@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                   �?���Q��?
             .@                                 �b@      �?              @                               ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �?��G���?-            �R@        ������������������������       �                     >@               &                   �`@�X����?             F@                                 �^@8�Z$���?             :@        ������������������������       �                     "@               %                    �?������?             1@                                    �?և���X�?             @        ������������������������       �                      @        !       "                   �_@���Q��?             @        ������������������������       �                      @        #       $                    @J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        '       2                    @X�<ݚ�?             2@       (       -                   `c@�n_Y�K�?
             *@       )       ,                 ����?�<ݚ�?             "@       *       +                    �M@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        .       /                   8p@      �?             @        ������������������������       �                      @        0       1                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�b��       h�h)h,K ��h.��R�(KK3KK��ha�B0  m��:m�?&�X�%�?�k(���?y�5���?UUUUUU�?UUUUUU�?              �?      �?        X|�W|��?���?J��yJ�?�־a��?W�+�ɕ?}g���Q�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?      �?                      �?�������?333333�?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?              �?#�u�)��?v�)�Y7�?      �?        �E]t��?]t�E]�?;�;��?;�;��?      �?        xxxxxx�?�?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?r�q��?;�;��?ى�؉��?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK'hyh)h,K ��h.��R�(KK'��h��B�	                             �?l�;�	�?[            �b@                     	             �?     ��?4             T@                                  �n@>���Rp�?             =@                                  �?j���� �?             1@        ������������������������       �                     @                                   �F@��
ц��?
             *@        ������������������������       �                     @               	                    �L@���Q��?             $@        ������������������������       �                     @        
                           @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@                                  �r@�IєX�?"            �I@                                  @`���i��?             F@       ������������������������       �                    �D@                                  �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?����X�?             @        ������������������������       �                     �?                                  �c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @               "       	             �?ףp=
�?'            �Q@                                  �?     �?$             P@                                    H@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                   c@0�)AU��?            �L@       ������������������������       �                    �H@                !                     L@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        #       $                   �l@�q�q�?             @        ������������������������       �                     @        %       &                    @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK'KK��ha�Bp  t�@�t�?ƒ_,���?      �?      �?GX�i���?�i��F�?ZZZZZZ�?�������?              �?�;�;�?�؉�؉�?      �?        �������?333333�?              �?�������?�������?      �?                      �?              �?�?�?F]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        �������?�������?      �?     ��?�$I�$I�?�m۶m��?      �?                      �?p�}��?��Gp�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhG        hNhEK
hGKhHh)h,K ��h.��R�(KK��ha�C              �?�t�bhThfhOC       ���R�hjKhkhnK
h)h,K ��h.��R�(KK��hO�C       �t�bK��R�}�(hKhxK/hyh)h,K ��h.��R�(KK/��h��B�                          pff�?���Q��?c            �b@                     	             �?ĴF���?4            �T@               
                    �?�q�q�?             (@                                  ^@      �?              @        ������������������������       �                     �?                                   @J@և���X�?             @        ������������������������       �                      @               	                   �k@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �g@hA� �?,            �Q@                                  �?0�,���?*            �P@                                 `a@0�)AU��?%            �L@       ������������������������       �                     D@                                   @N@�IєX�?
             1@       ������������������������       �        	             0@        ������������������������       �                     �?                                @33�?ףp=
�?             $@                                  @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                  pn@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               ,                   Xu@�M���?/             Q@              #                    �?��.��?-            �N@               "                   �c@���Q��?             $@              !                   �`@      �?              @                                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        $       '       	             �?�:�]��?%            �I@       %       &                   �e@�nkK�?!             G@       ������������������������       �                      F@        ������������������������       �                      @        (       +                    @���Q��?             @       )       *                 833@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        -       .                    �?����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK/KK��ha�B�  333333�?�������?E�JԮD�?ە�]�ڵ?UUUUUU�?UUUUUU�?      �?      �?              �?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?              �?        ���?_�_�?Ez�rv�?g��1��?��Gp�?p�}��?      �?        �?�?      �?                      �?�������?�������?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?<<<<<<�?�������?������?�����?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�?}}}}}}�?d!Y�B�?�Mozӛ�?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�m۶m��?�$I�$I�?      �?                      �?�t�bubhhubehhub.